
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka

include(lib_user.ckt);line 1.5; l_current(i_1,above,0.5); dot;       { line right_ 1 up_ 1; l_current(i_2,above rjust)};      line right_ 1 down_ 1;l_current(i_3,above ljust);
.PE
