.PS
scale=2.54
cct_init

include(base.ckt)
Grid(10,5);
move to (1,2);
bjt_NPN(1,1,L);
bjt_NPN(1,1,L,N);

bjt_PNP(1,1,L);
bjt_PNP(1,1,L,N);

move to (1,0.5);
bjt_NPN(1,1,R);
bjt_NPN(1,1,R,N);

bjt_PNP(1,1,R);
bjt_PNP(1,1,R,N);

move to (8, 1.25);
Q1: bjt_NPN(1.5, 1,L);
"\textit{Q1}" at Q1.e;
"\textit{Q1.B}" at Q1.B rjust;
"\textit{Q1.E}" at Q1.E below; 
"\textit{Q1.C}" at Q1.C above; 



.PE
