
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

#Grid(5,3.5);
Origin: Here 

box wid 2 ht 1 "Box";
line -> right_ 1;
circle rad 0.5 "r=0.5";
line -> right_ 1;
ellipse wid 2 ht 1 "Ellipse";


.PE
