
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)
Grid(8.5,2.5);
color_red;        # A. spline krivka, súradnic rovnake ako pri čiare
spline from (0,1.5) right_ 1 up_ 1 then right_ 0.5 down_ 1 then right_ 1 down_ 2 then up_ 3; "A" rjust below; 


color_blue;        # B. obojstranná šipka na krivke                       
spline <-> from (5.5,0) to (6,2) to (7,0.5) to (8.5,2); "B" rjust above; 


color_dark_green;  # C. Parameter tension
spline 1.4 from (3, 0.) up_ 2 then right_ 2 then down_ 2 dashed .08;
spline 1.0 from (3, 0.) up_ 2 then right_ 2 then down_ 2;
spline 0.6 from (3, 0.) up_ 2 then right_ 2 then down_ 2 dotted .05;"C" rjust above;

.PE
