
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


cct_init
log_init

include(lib_base.ckt)
include(lib_user.ckt)
include(lib_ic555.ckt)

command "\sf"

IC1: IC555_1 at (2,6.5); "555" at IC1.BX.n above;
IC2: IC555_2 at (7,6.5);
IC3: IC555_3 at (5,1);

.PE
