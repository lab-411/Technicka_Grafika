
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

Origin: Here 
move to (0.5, 1.5);   

resistor;           llabel(,R_1,); 
resistor(3,6,);     llabel(,R_2,); rlabel(,n=6,);  
resistor(,,Q);      llabel(,R_3,);   
resistor(,,H);      llabel(,R_4,); 

move to (0.5, 0.25); 

resistor(,,E);      llabel(,R_5,); 
resistor(,,ES);     llabel(,R_6,); 
resistor(,,V);      llabel(,R_7,); 
resistor(3,,E,1.5); llabel(,R_8,); rlabel(,linespec=3,);

.PE
