
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_color.ckt);
right_; 
resistor(2,,E); llabel(,R_1,); 

[  
      color_grey;
      boxrad=0.1
      box wid elen_ ht elen_*4/5 fill 0.95 ;
      color_reset;
      resistor(from last box.w to last box.e,, ES);
      llabel(,R_2,); rlabel(,470 \Omega / 5 W,);

]
resistor(2,,E); llabel(,R_3,);

.PE
