
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)
Grid(5,3);

    w=2;
    move to (1,1.5);                  # poloha zloženého objektu
A:[                                # blok s absolutnymi suradnicami  
        rr=0.25;                      # vnutorne premenne
        h=w/2; w=w+1/2;
    B:  box at (0,0) wid w ht h; 
    C1: circle at (0, 0.5) rad rr; 
    C2: circle at (0,-0.5) rad rr;
    C3: circle at B.w rad  rr;
    C4: circle at B.e rad rr;
] 

color_red;
r = A.C1.rad
line <- from A.B.nw left_ 1 up_ 1; "\sf A.B.nw" above;
line <- from A.ne right_ 1 up_ 1; "\sf A.ne" above;

right_; box at A.c wid A.wid_   ht A.ht_ dashed;

.PE
