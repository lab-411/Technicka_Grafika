
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)

Origin: Here 
Grid(10,5);


BOX: box wid 3 ht 2 at (5,3);
    "stred \,\,\,  boxu" at BOX.c;             dot;
    "\color{red} červený text" at BOX.n above; dot;

    color_dark_orange;
    "\color{blue} text vpravo" at BOX.e ljust; dot;
    "text vlavo dole" at BOX.sw rjust below;   dot;

    color_blue;
LL: line from (2, 0.5) right_ 6;
    "stred čiary" at last line.c above;        dot;

.PE
