
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


command"\sf"
include(lib_color.ckt)
include(lib_user.ckt)
include(lib_base.ckt)

right_;
move to (1,1.5);
T: d_fet(up_,,N);

color_red;
line <- from T.G left_ 0.75;    ".G" rjust;
line <- from T.D up_ 0.5 ;  ".D" above ;
line <- from T.S down_ 0.5;   ".S" below ;

right_;
color_black;
move to (4,1.5);


T: d_fet(up_,,P);
color_blue;
B: box wid (T.w-T.e).x ht (T.n-T.s).y at T.c dotted;
line <- from T.sw down_ 0.5 left_ 0.5;   ".sw" below rjust;
line <- from T.nw up_ 0.5 left_ 0.5;     ".nw" above rjust;
line <- from T.ne up_ 0.5 right_ 0.5;    ".ne" above ljust;
line <- from T.se down_ 0.5 right_ 0.5;  ".se" below ljust;
line <- from T.e  right_ 0.75;  ".e" ljust;
line <- from T.w  left_ 0.75;  ".w" rjust;
line <- from T.n  up_ 0.75;  ".n" above;
line <- from T.s  down_ 0.75;  ".s" below;
line <- from T.c  down_ 0.55 right_ 1.25;  ".c" ljust ;

.PE
