
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


resistor(2,,E); llabel(,\sf R_1,)
dot "\sf 3.3V" above; {resistor(down_ 2 ,,E);  llabel(,\sf R_3,)}
resistor(right_ 2,,E);  llabel(,\sf R_2,)

.PE
