
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


    include(lib_base.ckt)
    include(lib_color.ckt)
    #Grid(7,7);
    move to (4,2)
    up_;
T1: bi_tr(2, L, N,E); 
    resistor(from T1.E down_ 1.5,,E); rlabel(,R_e,);
GN: gnd;

RC: resistor(from T1.C up_ 1.5,,E); llabel(,R_c,);
DC: dot;
    tconn(0.75,O); clabel(,,V_+); 

    color_red
    line from T1.B left_ 0.8; 
D1: dot; dlabel(0,0,,V_b,,AL);
    resistor(from D1 down_ (D1.y - GN.n.y),,E); rlabel(,R_{b1},);
    gnd;
    color_black;

    resistor(from D1 up_ (RC.end.y - D1.y),,E); llabel(,R_{b2},); 
    line to DC;

    capacitor(from D1 left_ 1.5); rlabel(,C_{b},); 
    tconn(0.5,O); rlabel(,V_{in},);

    move to T1.C; 
D2: dot; dlabel(0,0,,V_c,,R);
    capacitor(from D2 right_ 1.5); llabel(,C_{c},); 
    tconn(0.5,O); llabel(,V_{out},);

    move to T1.E; 
D3: dot; dlabel(0,0,,V_e,,R); 
    line right_ 1;
    capacitor(down_ 1.5); llabel(,C_{e},); 
    gnd;

.PE
