
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


cct_init
log_init
include(lib_base.ckt)
include(lib_color.ckt)
include(lib_ic555.ckt)
command "\sf"
#Grid(6,6)

IC: IC555_2 at (3,3);
    C2: capacitor(from IC.Pin5 down_ 0.75,); llabel(,\sf 10nF,);
        line from IC.Pin7 left 1;
        dot;
        {R1: resistor(up_ 1.5,,E); llabel(,\sf R_1,); } #DT1: dot; }
        R2: resistor(down_ 1.5,,E); rlabel(,\sf R_2,); DT2: dot;
     C1: capacitor(1.25,); rlabel(,\sf C,); 
        line right_ to (IC.Pin1, Here); 
        dot;
        {line to IC.Pin1;}
        {line to (IC.Pin5, Here) then to C2.end; }
        down_; gnd(0.5);

    # vetva napajania
        line from R1.end to (IC.Pin4, R1.end);
        dot;
        {line to IC.Pin4;} 
        {line to (IC.Pin8, Here) then to IC.Pin8;}
        up_; power(0.75, $\sf V_{cc}$ );
    # vystup        
        move to IC.Pin3; right_; tconn(,O); "$\sf V_{out}$" at Here ljust;
        "555" at IC.BX.ne ljust below;

        d = (IC.Pin2.x - DT2.x)/2
        line from DT2 right_ d; line up_ to (Here, IC.Pin2); dot; 
        {line to IC.Pin2;} 
        line up_ to (Here, IC.Pin6) then to IC.Pin6;

.PE
