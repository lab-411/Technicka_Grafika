
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

Origin: Here 
move to (0.5, 1.5);   

capacitor;          llabel(,C_1,); 
capacitor(,C,);     llabel(,C_2,);    
capacitor(,E);      llabel(,C_3,); 
capacitor(,K);      llabel(,C_4,); 

move to (0.5, 0.0); 

capacitor(,M, ,0.75, 0.25);      llabel(,C_5,); 
capacitor(,P);      llabel(,C_6,);  
capacitor(, CP);    llabel(,C_7,);   
capacitor(,+LC);     llabel(,C_8,); 

.PE
