
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

Origin: Here 
Grid(3,3);
    right_;
    r = 1.5;
    move to (0,r);
C1: circle diam 2*r;
    color_red;
    alpha = pi_ / 4;     # uhol v radianoch
    line from C1.c to C1.c + (cos(alpha), sin(alpha))*r;
D1: dot;

.PE
