
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


    include(lib_base.ckt)
    Grid(15,5);
    move to (3,3);
OP: opamp()
    line from OP.In1 left 0.5;
DN: dot;
    resistor(2,,E); llabel(,R_1,);
    circle rad 0.1; "\textit{In}" at last circle.n above;

    line from DN up_ 1;
    resistor(right_ 2.5,,E); llabel(,R_2,);
    line down_ (Here.y - OP.Out.y);
DO: dot;
    { line to OP.Out; }
    line right_ 1;
    circle rad 0.1; "\textit{Out}" at last circle.n above;

    line from OP.In2 left_ 0.5 then down_ 0.5; gnd; 
    "\textit{Invertujúci zosilovač}" at OP.c + (0, -1.5);
    "$K = -\dfrac{R_2}{R_1}$" at OP.c + (0, -2.25);

move to OP.c + (6,0.5);
    right_;
PP: opamp(,,,,R)
    line from PP.In1 left_ 1.5;
    circle rad 0.1; "\textit{In}" at last circle.n above;
    line from PP.In2 left_ 0.5 then down_ 0.75;
    dot;
    {resistor(down_ 1.5,,E); rlabel(,R_1,); gnd;}
    resistor(right_ 2.5,,E); llabel(,R_2,);
    line up_ -(Here.y - PP.Out.y);
    dot;
    { line to PP.Out; }
    line right_ 1;
    circle rad 0.1; "\textit{Out}" at last circle.n above;
    "\textit{Neinvertujúci zosilovač}" at PP.c + (0, 1);
    "$K =1 + \dfrac{R_2}{R_1}$" at PP.c + (0.5, -2.25);

.PE
