.PS
scale = 2.54      
maxpswid = 30   
maxpsht = 30 
cct_init        

circle rad 1 fill 0.8
resistor();

.PE
