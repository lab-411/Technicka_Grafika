
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)
B1: box wid 2 ht 2;
line from B1.ne -(0,0.25) right_ 1 ;
P1: circle rad .1; "\textit{P1}" at P1.e ljust;

line from B1.se + (0,0.25) right_ 1 ;
P2: circle rad .1; "\textit{P2}" at P2.e ljust;

"\textit{Output}" at (P1 + P2)/2;

color_red;
"\small{ \"Output\" at (P1 + P2)/2;}" at B1.s + (0,-.2) below ljust;
line from B1.e + (.2, 0) right 2 dotted;
line from P1.s + (0, -0.1) to P2.n + (0,0.1) dotted;

.PE
