
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

Origin: Here 
move to (0.5, 1.5);   

diode;          llabel(,D_1,); 
diode(,S,);     llabel(,D_2,); rlabel(,S,);  
diode(,V);      llabel(,D_3,); rlabel(,V,);  
diode(,v);      llabel(,D_4,); rlabel(,v,);

move to (0.5, 0.25); 

diode(,U);     llabel(,D_5,); rlabel(,U,);  
diode(,ZK);    llabel(,D_6,); rlabel(,ZK,); 
diode(,T);     llabel(,D_7,); rlabel(,T,);  
diode(,,R);    llabel(,D_8,); rlabel(,Rev,);

.PE
