
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)
move to (3.5,0);

color_black; box wid 1 ht 0.5; "co\\lor\_black" at last box .w rjust;
color_grey; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_grey" at last box .w rjust;
color_blue; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_blue" at last box .w rjust;
color_green; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_green" at last box .w rjust;
color_red; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_red" at last box .w rjust;
color_olive; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_olive" at last box .w rjust;
color_khaki; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_khaki" at last box .w rjust;
color_dark_khaki; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_khaki" at last box .w rjust;
#color_lemonchiffon; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_lemonchiffon" at last box .w rjust;
color_steelblue; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_steelblue" at last box .w rjust;
#color_snow; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_snow" at last box .w rjust;
#color_honeydew; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_honeydew" at last box .w rjust;
#color_mintcream; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_mintcream" at last box .w rjust;

move to (5,0);

color_cyan; box wid 1 ht 0.5; "co\\lor\_cyan" at last box .e ljust;
color_brown; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_brown" at last box .e ljust;
color_orange; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_orange" at last box .e ljust;
color_violet; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_violet" at last box .e ljust;

color_light_grey; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_light\_grey" at last box .e ljust;
#color_light_yellow; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_light\_yellow" at last box .e ljust;
color_light_blue; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_light\_blue" at last box .e ljust;

color_dark_grey; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_grey" at last box .e ljust;
color_dark_cyan; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_cyan" at last box .e ljust;
color_dark_green; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_green" at last box .e ljust;
color_dark_orange; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_orange" at last box .e ljust;
color_dark_red; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_red" at last box .e ljust;
color_dark_violet; box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_dark\_violet" at last box .e ljust;

color_aquamarine;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_aquamarine" at last box .e ljust;
color_silver;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_silver" at last box .e ljust;
color_cadetblue;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_cadetblue" at last box .e ljust;
color_coral;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_coral" at last box .e ljust;
color_gold;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_gold" at last box .e ljust;
color_mediumForestGreen;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_mediumForestGreen" at last box .e ljust;
color_slategrey;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_slategrey" at last box .e ljust;
color_firebrick;  box wid 1 ht 0.5 with .ne at last box.se + (0, -0.1); "co\\lor\_firebrick" at last box .e ljust;

.PE
