
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

#Grid(6,1.5);
command "\sf"

ground(at (0.5,1),,N); "N" at last box above;
ground(at (1.5,1),,F); "F" at last box above;
ground(at (2.5,1),,S); "S" at last box above;
ground(at (3.5,1),,L); "L" at last box+(0,0.3) above;
ground(at (4.5,1),,P); "P" at last box+(0,0.3) above;
ground(at (5.5,1),,E,); "E" at last box above;

.PE
