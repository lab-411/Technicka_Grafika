      
.PS
cct_init               
                       
scale = 2.54           
maxpswid = 30          
maxpsht = 30           
arrowwid  = 0.127     
arrowht = 0.254        
boxrad = 0.1;
                        
include(lib_base.ckt)
include(lib_color.ckt)
include(lib_user.ckt)

Origin: Here 
command"\sf"

#move to (15, 10);

# TODO
# Doplnit napajacie zdroje
# doplnit znacky tenzometrov v mostiku
# doplnit oznacenie dynamometra
# doplnit CPU

#-----------------------------------------------------------------------
# Timer
#-----------------------------------------------------------------------
    down_;
ARR:box wid 4 ht 1; {"Auto-Reload Register" at last box.c;}
    line -> down_ 1;
    {
        LC: last line.c;
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "16" at LC + (-0.25 , 0) above;
    }

CC1:box wid 4 ht 1; {"Compare Register 1" at last box.c;}
    line -> from CC1.e right_ 3;
    {
        LC: last line.c + (0.5,0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "1" at LC + (-0.25 , 0) above;
            "pulse" at LC + (-0.25 , -0.55) above;
            move to LC + (-0.5, 0.75); {"$5 \mu s$" at Here + (0.35, 0.5) above;}
            line right_ 0.25 then up_ 0.5 then right_ 0.25 then down_ 0.5 then right_ .5;
    }

HB: box wid 2 ht 2; {"HBS57" at last box.c;}; # controller

    move to (ARR.w + CC1.w)/2 + (-0.5,0);
TIM:box wid 5 ht 3.5; {"TIM1" at last box.n above;}

    line <- from ARR.w left_ 1.5;
PRE:box wid 1 ht 1;  
    {
        ":N" at last box.c;
        "prescaler" at last box.n above;
    }
    line <- from last box.w left_ 1; "sysclk" at last line.end rjust;

#-----------------------------------------------------------------------
# Motor 
#-----------------------------------------------------------------------

    move to HB.n + (-0.75, 2);

MS: Here
    line up_ 0.5; right_; inductor(2,W,8); line down_ 0.5;
    move to MS + (-1,3); line right_ 0.5; down_; inductor(2,W,8);
    line left_ 0.5;
    move to MS + (2, 2);
MCC:circle rad 1;

    move to MCC.c; dot; # +(1.5/sqrt(2)/2, 0);
    Point_(45); rotbox(1.75, 0.25,thick 2, r=0.1) at MCC.c;

    move to MCC.c - (2, 0.25); right_;
MB: box wid 3.5 ht 3.5;                   # motor box
    {"stepper motor" at MB.n above;}

#-----------------------------------------------------------------------
# IRC
#-----------------------------------------------------------------------

    line -> from HB.n to MB.s;
    {
        LC: last line.c;
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "4" at LC + (-0.25 , 0) above;
    }

    line -> from MCC.c right_ 3.75 dashed invis;
    dot;
IRC:circle rad 1 with .c at last line.end; {"IRC" at IRC.n above;}

    #color_blue;
    for i=0 to pi_*2 by pi_/16 do  {line from (sin(i), cos(i) )*0.35 + IRC.c to (sin(i), cos(i) )*0.9 + IRC.c; }
    color_black;

    color_red;
    line -> from MCC.c to IRC.c dashed thick 1.5 ;
    color_black;

    line from IRC.s to (IRC.c.x, HB.e.y);
    {
        LC: last line.c;
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "4" at LC + (-0.25 , 0) above;
    }
    line -> to HB.e;

#-----------------------------------------------------------------------
# GPIO
#-----------------------------------------------------------------------

    move to TIM.s + (1.5, -1);
    down_;
GPIO:box wid 2 ht 1 ; {"GPIO" at last box.c;}
    line from GPIO.e to (HB.s.x, last box.c.y);
    {
        LC: last line.c;  # + (0.5, 0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "2" at LC + (-0.25 , 0) above;
            "direction, enable" at LC + (-0.25 , -0.55) above;
    }
    line -> to HB.s;

#-----------------------------------------------------------------------
# mostik a ADC prevodnik
#-----------------------------------------------------------------------

    move to PRE.c + (-6,3);
    right_; 
ADC: adc(2,1,2,,1,); 
    {   "24 bit" at ADC.c; 
        "ADC" at ADC.n + (0,0.1) above; 
        "MCP3651" at ADC.n + (0,0.45) above; 
    }

    line from ADC.In1 left_ 1.5; 

    DT1: dot;
    Point_(180-45) resistor(,E); 
    DT2: dot;
    Point_(180+45) resistor(,E);
    DT3: dot;
    Point_(-45) resistor(,E);
    DT4: dot;
    Point_(+45) resistor(,E);

    move to DT2; line up_ 0.25; power(0.5,3.3V);
    move to DT4; line down_ 0.25; gnd;

    line from ADC.In2 left_ 1 then down_ 2;
    line to (DT3.x - 0.5, Here.y);
    line to DT3-(0.5,0) then to DT3;

    line <-> from ADC.Out right_ 1.5;
    {
        LC: last line.c; # + (0.75,0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "4" at LC + (-0.25 , 0) above;
            box  at LC.c + (0,-.45)  wid 1 ht 0.45 "MISO" invis; down_;   
            box  wid 1 ht 0.45  "MOSI" with .n at last box.s invis;          
            box  wid 1 ht 0.45  "CLK" with .n at last box.s invis;
            box  wid 1 ht 0.45  "CS" with .n at last box.s invis;
    }

SPI: box wid 2 ht 1; {"SPI2" at last box.c;}
    move to SPI.e + (2,0);
RTC:box wid 2 ht 1; {"RTC" at last box.c;}

#-----------------------------------------------------------------------
# SDCARD
#-----------------------------------------------------------------------

    move to PRE.c + (-2.5,-4.25);
    right_;
SPI2: box wid 2 ht 1; {"SPI1" at last box.c;}
    line <-> from SPI2.w left_ 2; 
    {
        LC: last line.c; # + (0.75,0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "4" at LC + (-0.25 , 0) above;
            box  at LC.c + (0,-.45)  wid 1 ht 0.45 "MISO" invis; down_;   
            box  wid 1 ht 0.45  "MOSI" with .n at last box.s invis;          
            box  wid 1 ht 0.45  "CLK" with .n at last box.s invis;
            box  wid 1 ht 0.45  "CS" with .n at last box.s invis;
    }

    dcx = 0.2;    # sdkarta
    dch = 0.5;
    dcl = 1.7
    line up dch;
    line to Here+ (-dcx, dcx);
    line left dcl;
    line down (dch+dcx)*2 then right dcl+dcx;
    line up dch+dcx;
    {"SDCARD" at Here - ((dcl+dcx)/2, 0);}



#box wid 2 ht 1; 
# {
#    "Display" at last box.c above;
#    "Keyboard" at last box.c below;
# }

#-----------------------------------------------------------------------
# USART
#-----------------------------------------------------------------------
    move to PRE.c + (-2.5,-2.25);
    right_;
USART: box wid 2 ht 1;
    {"USART2" at last box.c;}
    line <-> from USART.w left_ 2; 
    {
        LC: last line.c; # + (0.75,0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "2" at LC + (-0.25 , 0) above;
            "Rx" at LC.c + (0, -0.55) above;
            "Tx" at LC.c + (0, -0.95) above;
    }
    box wid 1 ht 1; 
    line from last box.sw to last box.ne; {"USB / TTL" at last box.n above;}
    line -> from last box.w left_ 2; {"USB" at last line.end rjust;}

#-----------------------------------------------------------------------
# Koncove spinace
#-----------------------------------------------------------------------
    line <- from GPIO.s  down_ 1.5;
    line to (HB.w.x, Here.y);
    {
        LC: last line.c + (0.75,0);
            line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
            "2" at LC + (-0.25 , 0) above;
            "swi\\tch" at LC + (-0.25 , -0.55) above;
    }
    right_;
    box wid 2 ht 2; 
    move to last box.w + (0, 0.5); single_switch(2, OFF, H);
    move to last box.w + (0, -0.5); single_switch(2, OFF, H);

#-----------------------------------------------------------------------
# SPI periferie
#-----------------------------------------------------------------------

    move to PRE.c + (-2.5,-6.25);
    right_;
I2C: box wid 2 ht 1; {"I2C1" at last box.c;}
    line <- from I2C.s down 1.5;

    {
        LC: last line.c #  + (0.75,0);
         line from LC-(0.15, 0.15) to LC+(0.15, 0.15)
         "2" at LC + (-0.25 , 0) above;
         "SCK, SDL" at LC + (+0.2 , 0.0) ljust;
    }

DT1:dot;
    {
            line -> left 3 then down 0.5;
      KEYB: box wid 1.5 ht 1;
            "KEYB" at last box.c;
    }

    {
            move from DT1 left 1;
            line -> down 0.5;
        DISP: box wid 1.5 ht 1;
            "DISP" at last box.c;
    }

    {
        line -> right 3 then down 0.5;
      LEDS: box wid 1.5 ht 1;
        "LEDS" at last box.c;
    }

    {
            move from DT1 right 1;
            line -> down 0.5;
        TEMP: box wid 1.5 ht 1;
            "TEMP" at last box.c;
    }

#-----------------------------------------------------------------------
# ramik
#-----------------------------------------------------------------------
    bw = 9+1/2;
    bh = 10+3/4;

    move to (SPI.nw)+ (-1/4, -bh/2+1/4);
    right_;
    color_red;
    boxrad = 0.25;
    box wid bw ht bh dashed thick 0.35;  {"STM32L476" at last box.n above;}
    color_black;
.PE
