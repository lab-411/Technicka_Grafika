
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)
Grid(4,4)

define(`triangle', `
[  
    line from (1,1) to (0,0) then to (1,-1);
    arc cw from (1,1) to (1,-1)
]')

move to (1,2);
color_red;
rgbfill(fill_yellow, {triangle} );

.PE
