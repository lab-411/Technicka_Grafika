.PS
scale=2.54
cct_init
include(base.ckt)
Grid(11.5,4);

# Usual defs...
move to (.6,3);
qrt=2;
hlf=0.5;

Q1:e_fet(up_ ,,,);   
move right_ hlf
Q2:e_fet(up_ ,R); 
move right_ hlf
Q3:e_fet(up_,,P)
move right_ hlf
Q4:e_fet(up_,R,P); 

move right_ hlf
Q5:d_fet(up_)
move right_ hlf
Q6:d_fet(up_,R)
move right_ hlf
Q7:d_fet(up_,,P)
move right_ hlf
Q8:d_fet(up_,R,P)
 
move to (0.35,1);
e_fet(up_,,,S)
move right_ hlf
e_fet(up_,R,,S)
move right_ hlf
e_fet(up_,,P,S)
move right_ hlf
e_fet(up_,R,P,S)
move right_ hlf
d_fet(up_,,,S)
move right_ hlf
d_fet(up_,R,,S)
move right_ hlf
d_fet(up_,,P,S)
move right_ hlf
d_fet(up_,R,P,S)

.PE
