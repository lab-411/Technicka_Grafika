
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_color.ckt)
include(lib_base.ckt)
Grid(5,3)

"\fbox{\color{red} Text v rámiku}" at (2.5, 0.5)

color_blue;
"\fbox{\large Text large v rámiku}" at (2.5, 1.5)

color_reset;
"\sf \fbox{\Large Text {\color{red} Large} v rámiku}" at (2.5 ,2.5)

.PE
