
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka



include(lib_base.ckt)
include(lib_user.ckt)
include(lib_color.ckt)

     move to (3,1);
T2:  bjt_PNP(0.6,1,R,N); {"$T2$" at T2.c + (-0.4, 0.5);}

     line from T2.E right 0.8; 
T22: bjt_PNP(1,1,R,N);    {"$T22$" at T22.e;}
     resistor(from T22.E left_ (T22.E.x - T2.E.x),,E); {rlabel(,R_2,);}
     line to T2.E; dot;

     line from T2.C right_ -(Here.x - T22.C.x); 
     dot; {line -> down_ 0.8;  "V-" below; }
     line to T22.C;

     move to T22.E; dot;
     line up_ 0.8; 
     dot; {line right_ 1.5; C1: circle rad 0.1}
     line up_ 0.8; 
     color_red;
DV:  dot;   { line <- from Here+(.1,0) to Here+(1,0); "DV" at Here ljust; }


T11: bjt_NPN(1,1,R,N) with .E at Here;     {"$T11$" at T11.e;}
     line from T11.B left_ 0.8;
T1:  bjt_NPN(0.6,1,R,N) with .E at Here;  {"$T1$" at T1.c + (-0.4, 0.5);}
     resistor(from T11.E left_ (T11.E.x - T1.E.x),,E); {llabel(,R_1,);} 
     line to T1.E; dot;
     color_black;

     line from T1.C right_ -(Here.x - T11.C.x); 
     dot; {line -> up_ 0.8;  "V+" above; }
     line to T11.C

     move to T1.B;
     down_;
DC:  dc_source( (T1.B.y - C1.c.y), 0.8, P); { line <- from DC.C.c+(-0.5,-0.5) to DC.C.c+(-0.5,0.5) "$V_1$" rjust}
     dot; {line left_ 1.5; C2: circle rad 0.1;}
     line to T2.B;

     line -> from C1.c + (0, -0.2) down_ 1 "$V_{out}$" ljust; circle rad 0.1 at Here + (0, -0.2); line down_ 0.25; gnd;
     line -> from C2.c + (0, -0.2) down_ 1 "$V_{in}$" ljust; circle rad 0.1 at Here + (0, -0.2); line down_ 0.25; gnd;

.PE
