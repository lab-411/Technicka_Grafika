
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_user.ckt)
command"\sf"
#Grid(10, 2.5);

move to (0.5, 2);
Q1:bjt_NPN(1,1,L);   {"Q1" at Q1.n above; }
Q2:bjt_NPN(1,1,L,N); {"Q2" at Q2.n above; }

Q3:bjt_PNP(1,1,L);   {"Q3" at Q3.n above; }
Q4:bjt_PNP(1,1,L,N); {"Q4" at Q4.n above; }

move to (0.5, 0.5);
Q5:bjt_NPN(1,1,R);   {"Q5" at Q5.s below; }
Q6:bjt_NPN(1,1,R,N); {"Q6" at Q6.s below; }

Q7:bjt_PNP(1,1,R);   {"Q7" at Q7.s below; }
Q8:bjt_PNP(1,1,R,N); {"Q8" at Q8.s below; }

move to (9, 1.25);
Q10: bjt_NPN(1.5, 1, R);
"\textit{Q10}" at Q10.e;
"\textit{Q10.B}" at Q10.B rjust;
"\textit{Q10.E}" at Q10.E below; 
"\textit{Q10.C}" at Q10.C above; 

.PE
