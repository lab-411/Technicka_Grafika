define(`IC485', `[
  BX: box wid 2 ht 5*lg_pinsep;

      lg_pin(BX.nw - (0, 1*lg_pinsep), RO, Pin1, w, 1);
      lg_pin(BX.nw - (0, 2*lg_pinsep), lg_bartxt(RE), Pin2, wN, 2);
      lg_pin(BX.nw - (0, 3*lg_pinsep), DE, Pin3, w, 3);
      lg_pin(BX.nw - (0, 4*lg_pinsep), DI, Pin4, w, 4);

      lg_pin(BX.ne - (0, 1*lg_pinsep),  Vcc, Pin8, e, 8);
      lg_pin(BX.ne - (0, 2*lg_pinsep),  lg_bartxt(B), Pin7, eN, 7);
      lg_pin(BX.ne - (0, 3*lg_pinsep),  A, Pin6, e, 6);
      lg_pin(BX.ne - (0, 4*lg_pinsep),  GND, Pin6, e, 5);
      
      arc ccw from BX.n-(.2,0) to BX.n+(0.2,0) with .c at BX.n;
      rgbfill(fill_black, {circle at BX.nw + (0.15, -0.15) rad 0.055} )
]')

define(`IC485_LEFT', `[
  P1: (-1.5,  1.00);
  P2: (-1.5,  0.33);
  P3: (-1.5, -0.33);
  P4: (-1.5, -1.00);
  P7: ( 0.5,  0.33);
  P6: ( 0.5, -0.33);
  
    rgbfill(fill_light_yellow, { BX: box wid 2 ht 3.25 at (-0.5,0);})
    lg_pin( P1,,Pin1,w,RO);
    lg_pin( P2,,Pin2,w,lg_bartxt(RE));
    lg_pin( P3,,Pin3,w,DE);
    lg_pin( P4,,Pin4,w,DI);
    lg_pin( P7,,Pin7,e,lg_bartxt(B));
    lg_pin( P6,,Pin6,e,A);
  
    color_red;
    left_
  BR:  BUFFER_gen(TOC, 0.9, 0.9,NP,N,,, ) with .Out at P1+(0.25,0); "R" at BR.C;
    right_
  BD: BUFFER_gen(TC,0.9, 0.9,P,PN,P,,) with .In1 at P4+(0.3,0); "D" at BD.C;
    color_black;
    line from BD.SE1 right_ 1;  line to (Here, P3);
  DT1: dot; line to (Here, BR.In2) then to BR.In2
    line from BD.NE2 -(-0.05, 0.08) right_ 0.35; line to (Here, P2);
  DT2: dot; line to (Here, BR.In1) then to BR.In1
    line from BD.NE1 to (BD.NE1, P3) then to P3;
    line from BR.N_NE1 + (0, -0.05)to (BR.N_NE1 , P2) then to P2;
    line from BR.Out to P1;
    line from BD.In1 to P4;
    line from DT1 to P6;
    line from DT2 to P7;
]')


define(`IC485_RIGHT', `[
  P1: ( 1.5,  -1.00);
  P2: ( 1.5,  -0.33);
  P3: ( 1.5,  0.33);
  P4: ( 1.5,  1.00);
  P7: (-0.5,  0.33);
  P6: (-0.5,  -0.33);
  
    rgbfill(fill_light_yellow, { BX: box wid 2 ht 3.25 at (0.5,0);})
    lg_pin( P1,,Pin1,e,RO);
    lg_pin( P2,,Pin2,e,lg_bartxt(RE));
    lg_pin( P3,,Pin3,e,DE);
    lg_pin( P4,,Pin4,e,DI);
    lg_pin( P7,,Pin7,w,lg_bartxt(B));
    lg_pin( P6,,Pin6,w,A);
   
    color_red;
    right_
  BR:  BUFFER_gen(TOC, 0.9, 0.9,NP,N,,, ) with .Out at P1+(-0.25,0); "R" at BR.C;
    left_
  BD: BUFFER_gen(TC,0.9, 0.9,P,PN,P,,) with .In1 at P4+(-0.3,0); "D" at BD.C;
    color_black;
     line from BD.SE1 left_ 1;  line to (Here, P6);
  DT1: dot; line to (Here, BR.In2) then to BR.In2;

    line from BD.NE2 +(-0.05, 0.08) left_ 0.35; line to (Here, P7);
  DT2: dot; line to (Here, BR.In1) then to BR.In1;
    line from BD.NE1 to (BD.NE1, P3) then to P3;
    line from BR.N_NE1 + (0, 0.05)to (BR.N_NE1 , P2) then to P2;
    line from BR.Out to P1;
    line from BD.In1 to P4;
    line from DT1 to P6;
    line from DT2 to P7;
]')


define(`LINE_485', `[
  spline 1.0 from (0, 0.33)   to (0.5, 0.33) to (1., -0.43) to (1.5, 0.43) to (2., -0.43) to (2.5, 0.33) to (3, 0.33);
  spline 1.0 from (0, -0.33)  to (0.5, -0.33) to (1., 0.43) to (1.5, -0.43) to (2., 0.43) to (2.5, -0.33) to (3, -0.33);
]')


define(`TERM_485', `[
    line from (0, 0.33) right_ 0.1;
    dot;
    {line right_ 1.5;}
    line down_ 0.33; resistor(right_ 1.3,,E); line down_ 0.33
    line from (0, -0.33) right_ 1.4; dot; line 0.2;
  ]')


