
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
"tb\\ox()" at (1.5, 3);
"tc\\onn()" at (4, 3);

move to (0.5,1.0); line 1; tbox(V_1, 1, , <); 
move to (0.5,1.5); tbox(V_2, 1, , >); line 1
move to (0.5,2.0); line 1; tbox(V_3, 1, , <>, fill_(0.9))

move to (3.5,0.5); T1: tconn(,O); "$0$" at T1.e ljust
move to (3.5,1.0); T2: tconn(,>); "$>$" at T2.e ljust
move to (3.5,1.5); T3: tconn(,<); "$<$" at T3.e ljust
move to (3.5,2.0); T4: tconn(,A); "$A$" at T4.e ljust
move to (3.5,2.5); T5: tconn(,M); "$M$" at T5.e ljust

.PE
