
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

Origin: Here 
d = 2;
move to (2, 3);
DT1: dot;                   # referencny bod
{
         diode(right_ up_); dlabel(0,0,,D_1,,XAR);
    DT2: dot;              
         diode(right_ down_); dlabel(0,0,,D_2,,XAL);
}

{
         diode(right_ down_);   dlabel(0,0,,D_3,,XBR);
    DT3: dot;
         diode(right_ up_);    dlabel(0,0,,D_4,,XBL);
    DT4: dot;
}

# pouzitie referencii vytvorenych v blokoch
L1: line from DT2  up_ d/2 then left_ d;   tconn(,O);
L2: line from DT3  down_ d/2 then left_ d; tconn(,O);
L3: line from DT4 right_ d; tconn(d/4, O);
L4: line from DT1 left_ d/2 then down_ 7*d/8; 
    line to (L3.e.x, Here.y); tconn(right_ d/4,O);

.PE
