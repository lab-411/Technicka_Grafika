
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_user.ckt)

Grid(12,2);
move to (.5,1);
hlf=0.5;

Q1:bi_tr(up_ );   
move right_ hlf
Q2:bi_tr(up_ ,R); 
move right_ hlf
Q3:bi_tr(up_,,,E)
move right_ hlf
Q4:bi_tr(up_,R,,E); 

move right_ hlf
Q5:bi_tr(up_,,P)
move right_ hlf
Q6:bi_tr(up_,R,P)
move right_ hlf
Q7:bi_tr(up_,,P,E)
move right_ hlf
Q8:bi_tr(up_,R,P,E)

.PE
