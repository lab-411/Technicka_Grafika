
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


cct_init
log_init
include(lib_base.ckt)
include(lib_color.ckt)
include(lib_ic555.ckt)
command "\sf"

IC: IC555_2;
    line from IC.Pin7 left 1;
    dot;
    {R1: resistor(up_ 1.5,,E); llabel(,\sf R_1,); DT1: dot; }
     R2: resistor(down_ 1.5,,E); rlabel(,\sf R_2,); DT2: dot;
     C1: capacitor(1,); rlabel(,\sf C,); gnd();


     move to IC.Pin5; C2: capacitor(0.75,); llabel(,\sf 10nF,); gnd();
     move to IC.Pin1; gnd(0.5);

.PE
