.PS
scale=2.54
cct_init

include(base.ckt)
Grid(4,4)


define(`triangle', `
[  
    line from (1,1) to (0,0) then to (1,-1);
    arc cw from (1,1) to (1,-1)
]')

move to 1,2
color_red;
rgbfill(fill_yellow, {triangle} );


.PE
