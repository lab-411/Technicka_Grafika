
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
Origin: Here 

B: box wid 4 ht 2 

move to B.west;   "B.w"  rjust;    # rovnako ako B.w
move to B.c;      "B.c";    
move to B.e;      "B.e"  ljust;   
move to B.n;      "B.n"  above; 
move to B.s;      "B.s"  below;

move to B.ne;     "B.ne"  above ljust; 
move to B.nw;     "B.nw"  above rjust; 

move to B.se;     "B.se"  below ljust; 
move to B.sw;     "B.sw"  below rjust; 

.PE
