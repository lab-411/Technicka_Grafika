
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


command "\sf"
up_
Orig: Here
source ; dlabel(1.3,0,"( )")
move to (Orig+(1,0)); source(,AC,,,); dlabel(1.3,0,"AC")
move to (Orig+(2,0)); source(,G,,,); dlabel(1.3,0,"G")
move to (Orig+(3,0)); source(,H,,,); dlabel(1.3,0,"H")
move to (Orig+(4,0)); source(,I,,,); dlabel(1.3,0,"I")
move to (Orig+(5,0)); source(,P,,,); dlabel(1.3,0,"P")
move to (Orig+(6,0)); source(,R,,,); dlabel(1.3,0,"R")
move to (Orig+(7,0)); source(,T,,,); dlabel(1.3,0,"T")
move to (Orig+(8,0)); source(,U,,,); dlabel(1.3,0,"U")

.PE
