
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)
Grid(5,3);

move to (1, 1.5);

A:[  # absolutne suradnice v bloku 
    B: box at (0,0) wid 2 ht 1; 
   C1: circle at (0, 0.5) rad 0.25; 
   C2: circle at (0,-0.5) rad 0.25;
   C3: circle at B.w rad 0.25;
   C4: circle at B.e rad 0.25;
  ]

color_red;
box at A.c wid A.wid_ ht A.ht_ dashed;  # outer contour

.PE
