
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)
Grid(11.5,4);

# Usual defs...
move to (.6,3);
hlf=0.5;

Q1:e_fet(up_ ,,P,S);   
move right_ hlf
Q2:e_fet(up_ ,R); 
move right_ hlf
Q3:e_fet(up_,,P)
move right_ hlf
Q4:e_fet(up_,R,P); 

move right_ hlf
Q5:d_fet(up_)
move right_ hlf
Q6:d_fet(up_,R)
move right_ hlf
Q7:d_fet(up_,,P)
move right_ hlf
Q8:d_fet(up_,R,P)

move to (0.35,1);
e_fet(up_,,,S)
move right_ hlf
e_fet(up_,R,,S)
move right_ hlf
e_fet(up_,,P,S)
move right_ hlf
e_fet(up_,R,P,S)
move right_ hlf
d_fet(up_,,,S)
move right_ hlf
d_fet(up_,R,,S)
move right_ hlf
d_fet(up_,,P,S)
move right_ hlf
d_fet(up_,R,P,S)

.PE
