
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

Origin: Here 
move to (0.5, 1.5);   

inductor;          llabel(,L_1,); dot;
inductor(,W);      llabel(,L_2,); rlabel(,W,);  dot;  
inductor(,L);      llabel(,L_3,); rlabel(,L,);  dot;
L4: inductor(,L,6);     llabel(,L_4,); "L,6" at L4.center + (0,-.05) below;  

.PE
