
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
cct_init
log_init

define(`IN3', `
   line left_ 0.25 from $1.In1;
   line left_ 0.25 from $1.In2;
   line left_ 0.25 from $1.In3;
   line right_ 0.25 from $1.Out;
   move to last line.end + (0.5,0)
')

define(`IN2', `
   line left_ 0.25 from $1.In1;
   line left_ 0.25 from $1.In2;
   line right_ 0.25 from $1.Out;
   move to last line.end + (0.5,0)
')

# Enter your drawing code here
right_;
G1: AND_gate(3); IN3(G1);
G2: NAND_gate(3); IN3(G2);
G3: OR_gate(2); IN2(G3);
G4: NOR_gate(3); IN3(G4);
G5: NXOR_gate(2); IN2(G5);
#G6: NOT_gate(2,,0.8,0.8); line from G6.In1 up_ 1;

define(`conn', `
    line from $1 left_ (($1 - $2)/2).x;
    line up_ to (Here.x, $2.y) then to $2;
')


G1: AND_gate(2) at (5, 2); "\sf G1" at G1.n above;
G2: AND_gate(2) at (5, 0.5); "\sf G2" at G2.n above;
G3: OR_gate(2) at (7, (G1.c.y + G2.c.y)/2 ); "\sf G3" at G3.n above;
G4: NOT_gate() at (3.5, 2.5); "\sf G4" at G4.n above;
    conn(G3.In1, G1.Out)
    conn(G3.In2, G2.Out)
    conn(G1.In1, G4.Out)

    line from G4.In1 left_ 0.35; DT: dot; line left_ 0.5; "\sf Q" at last line.end rjust;
    line from G1.In2 to (LL.end.x, G1.In2.y); "\sf D1" at last line.end rjust; 
    line from G2.In2 to (LL.end.x, G2.In2.y); "\sf D0" at last line.end rjust;  
    line from G2.In1 to (DT.x, G2.In1.y) then to DT;
    line from G3.Out right_ 1;  "\sf Y" at last line.end ljust;

.PE
