.PS
scale=2.54
cct_init

include(base.ckt)
Grid(10,5);
up_
    move to (2,0)
    gnd;
SW: single_switch(2, OFF, V, L);
    dot; {line -> right 2; "\sf PC13" at last line .end ljust}
    resistor(1.5, ,E);
    power($\sf V_{dd}$)
    "\sf Blue Button" at SW.e ljust
    
move to (6,0);
gnd;
DD: diode(2,,R); { em_arrows(,-45, .35) at DD.center +(.3,-.3); }
    dot; {line -> right 2; "\sf PA5" at last line .end ljust}
    resistor(1.5, ,E);
    power($\sf V_{dd}$)
    "\sf Green LED" at DD.center + (.5,0) ljust 
   

.PE
