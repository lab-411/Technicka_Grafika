.PS
scale=2.54
cct_init
command"\small \sf"
include(lib_color.ckt)


move to (0,0); 
right_;
color_black();
OP: opamp(,,,,R);
# color_grey();
#box wid (OP.ne-OP.nw).x ht (OP.nw-OP.sw).y at OP.c dashed;
#color_blue();

line from OP.In1 left_ 0.5;# "2" above;
line from OP.In2 left_ 0.5; #"3" above;
P1: 0.25 between OP.N and OP.E;
P8:  0.5 between OP.N and OP.E;

P5: 0.75 between OP.S and OP.E;
#P4: 1/3 between OP.S and OP.E;
#P6: 2/3 between OP.S and OP.E;

line from P1 up_ 0.25;
line from P8 up_ 0.25;

C1: circle rad 0.095 with .n at P5+(0,-0.035) 
#line from P5 up_ 0.25;

#line from P4 down_ 0.25;
#line from P6 down_ 0.25;

.PE
