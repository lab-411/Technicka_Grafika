
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

TR: transformer(down_ 2,L,7,W,4);
"1" at TR.P1 rjust below;
"2" at TR.P2 rjust above;
"3" at TR.S1 ljust above;
"4" at TR.S2 ljust below;
"$TR_1$" at TR.n above;

line from TR.P1 left_ 1; 
TC1: tconn(0.5,O);
line from TR.P2 left_ 1; 
TC2: tconn(0.5,O);

line from TR.S1 up_ to (TR.S1.x, TC1.y) then right_ 0.5;
D1: diode(1); llabel(,D_1,) 
DT1: dot;
{tconn(1, O); }
{C1: capacitor(down_ 2); llabel(,C_1,) }
line from TR.S2 down_ to (TR.S2.x, TC2.y) then to C1.end;
DT2: dot;
{tconn(right_ 1, O); }

.PE
