.PS
scale=2.54
cct_init

include(base.ckt)
#Grid(10,10);
move to (2,2);

T3: bjt_NPN(0.6, 1, L, N); {"$T_3$" at T3.w ljust};  dot;
T4: bjt_NPN(0.6, 1, R, N); {"$T_4$" at T4.e rjust};

resistor(down_ 1.5 from T3.E,,E); rlabel(,1k,); line -> down_ 0.5; "$-$" at last line.end  below rjust
resistor(down_ 1.5 from T4.E,,E); llabel(,1k,); line -> down_ 0.5; "$-$" at last line.end  below rjust

# kolektory vstupn0ho dielu
move to T3.C; 
line up_ 0.75; 
Q3: dot; {line to (T3.B, Here) then to T3.B;}
line up_ 2;
T1: bjt_PNP(0.6, 1, R, N) with .C at Here; "$T_1$" at T1.e rjust;

move to T4.C; 
line to (Here, Q3); 
Q4: dot;
line up_ to (Here, T1.C);
T2: bjt_PNP(0.6, 1, L, N) with .C at Here; "$T_2$" at T2.w ljust;

line  from T1.E right_ (T2.E.x - T1.E.x)/2; dot; 
{reversed(`source',up_ 2,I); llabel(,I_k = 20 \mu A,);line -> up_ 0.5; "$+$" at last line.end ljust; }
line to T2.E;

# vstupne terminaly
line from T1.B left_ 0.5;
C1: circle rad 0.1;
 line -> from C1.c + (0, -0.2) down_ 0.75 "$U_{N}$" ljust; circle rad 0.1 at Here + (0, -0.2); line down_ 0.25; gnd;

line from T2.B right_ 0.5;
C2: circle rad 0.1;
 line -> from C2.c + (0, -0.2) down_ 0.75 "$U_{P}$" ljust; circle rad 0.1 at Here + (0, -0.2); line down_ 0.25; gnd;

# koncovy stupen
line from Q4 right_ 2.5; b_current("$I_1$",below_,,E,1);
QQ: dot; line 0.15;

T5: bjt_NPN(.6,1,R,N);  {"$T_5$" at T5.e rjust};
line from T5.E right_ 0.05;
T6: bjt_NPN(.6,1,R,N);  {"$T_6$" at T6.e rjust};
line -> from T6.E down_ 1; "$-$" at last line.end  below rjust
line from T5.C to (T6.C, T5.C); dot; {line to T6.C;}
line up_ 1;
Q5: dot; {diode(up_ 0.5, ,R); diode(up_ 0.5, ,R); DD: dot;}
line right_ 0.5; 
T8: bjt_PNP(1,1,R,N); move to T8.E; dot; line right_ 1; C3: circle rad 0.1;
    line -> from C3.c + (0, -0.2) down_ 0.75 "$U_{a}$" ljust; circle rad 0.1 at Here + (0, -0.2); line down_ 0.25; gnd;
T9: bjt_NPN(1,1,R,N) with .E at T8.E; line from T9.B to DD;

LA: line from Q5 left_ 0.95 dashed;
LB: line from QQ up_ to (QQ,Q5) then right_ 0.95 dashed;
CC: capacitor(from LA.end to LB.end ); llabel(,C_k,); rlabel(,30pF,)

# napajanie koncoveho stupna
line -> from T8.C down_ 0.75; "$-$" at last line.end rjust;
line -> from T9.C up_   0.75; "$+$" at last line.end rjust;
move to DD;
{reversed(`source',up_ 2,I); llabel(,I_2 = 300 \mu A,);line -> up_ 0.5; "$+$" at last line.end ljust; }
.PE
