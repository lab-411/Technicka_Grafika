.PS
scale=2.54
cct_init

l=elen_
# Enter your drawing code here
# \graphicspath{ {/home/pf/ownCloud/Share-Projekty/1010_GitHub_lab-411/Technicka_Grafika/
"\graphicspath{ {/home/pf/ownCloud/Share-Projekty/1010_GitHub_lab-411/Technicka_Grafika/src} } \includegraphics{cm_0905c.png}" at (1,1);


.PE
