
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
Grid(10.5,5);


"\textit{Italic 123}" at (1.5, 0.5);
"\textbf{Bold 123}" at (1.5, 1.0);
"\textsc{SmallCaps 123}" at (1.5, 1.5);
"\textsl{Slanted 123}" at (1.5, 2);
"\textrm{Roman 123}" at (1.5, 3.5);
"\textsf{Sans Serif 123}" at (1.5, 4);
"\texttt{Typewriter 123}" at (1.5, 4.5);

for i=0 to 300 by 60 do {
  move to ( 5 + 1*cos(i/180*pi), 2.5 + 1*sin(i/180*pi) );
  sprintf("\rotatebox{%g}{Text %g}", i,i );
}

"\tiny  tiny  \scriptsize scriptsize \footnotesize footnotesize" at (8.5, 4.5);
" \small small \normalsize normalsize " at (8.5,4)
"\large large  \Large Large " at (8.5,3.25)
"\LARGE LARGE" at (8.5,2.5)
"\huge huge" at (8.5, 1.5)
"\Huge Huge" at (8.5, 0.5)

.PE
