
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
include(lib_color.ckt)
define(`xc', `
  {
   Q: Here; line from Q+(-.1,-.1) to Q+(0.1, 0.1); 
   line from Q+(-.1, .1) to Q+(0.1, -0.1);
   circle at Q rad 0.1*1.4; 
   color_black;
   }
')

Grid(7,3);

circle at (0.5,2.5)rad 0.25 "1"
right_; move to (1,2.5); color_red; xc;
resistor(2);    # (1)

circle at (0.5,1.5)rad 0.25 "2"
move to (2,1.5); color_red; xc;
resistor(at (2,1.5) right_ 2,,E)


circle at (0.5, 0.5)rad 0.25 "3";
move to (1,0.5); color_red; xc;
resistor(right_ 2 from (1,0.5))

circle at (6.5, 2.5)rad 0.25 "4"; move to (6,2.5); color_red; xc;
move to (4,2.5); color_blue; xc;
RA: resistor(right_ 2); llabel(,R_a,); 
RB: resistor(down_ 2); llabel(,R_b,); color_blue; xc;
resistor(from RA.start to RB.end)
circle at (4.65, 1.15)rad 0.25 "5"; 

.PE
