
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

command "\sf"
gnd(0.5,D); move to Here +(0.5,0)
gnd(0.5, L); move to Here +(0.5,0)
gnd(0.5, R); move to Here +(0.5,0)
gnd(0.5, U); move to Here +(0.5,0)

power(0.75, Vcc, U);move to Here +(0.5,0)
power(0.75, Vcc, D);move to Here +(1,0)
power(0.75, Vcc, L);move to Here +(0.5,0)
power(0.75, Vcc, R);move to Here +(0.75,0)

.PE
