.PS
scale=2.54
cct_init


include(base.ckt)
Grid(6,7);


#-----------------------------------------------------------------------
# NPN - bipolárny tranzistor
# bjt_NPN(length_ce, length_b, L|R|U|D)
# length_ce   - dlzka vyvodov medzi C a E
# length_b    - dlzka vyvodu b
# L|R|U|D     - orientacia, todo U|D
#-----------------------------------------------------------------------
define(`bjt_NPN',`[

    ifelse(defn(`d'),  $1, d=1,  d=$1)     # dlzka CE
    ifelse(defn(`bx'), $2, bx=1, bx=$2)    # dlzka bazy
    
    define(dir, index(`RLUP',$3, 0) )    
    Q:box ht d wid 1.5 dotted #invis;
    dx = 0.5
    dv = 0.3;

    ifelse( eval(dir), 0, {
        CC: Q.w  + (0.5,0);
            x = linethick;
            linethick = 2;
            line from CC + (0.025, 0) up_ .20;
            line from CC + (0.025, 0) down_ .20;
            linethick = x;

            line from CC to CC + (0.5, dv)  then to CC + (0.5,  d/2);
            line from CC to CC + (0.5,-dv)  then to CC + (0.5, -d/2);
            line from CC to CC + (0.5-bx, 0);    # vyvod bazy

            dr = sqrt((0.5*0.5) + (dv*dv))
            pd = asin(dv/dr);
            dp = 20
            ph = pi - pd + pi/dp

            sy = 0.25*sin(ph) -dv
            sx = 0.25*cos(ph) +0.5
            line from CC + (0.5, -dv) to CC + (sx, sy); round;

            ph = pi - pd - pi/dp
            sy = 0.25*sin(ph) -dv
            sx = 0.25*cos(ph) + 0.5
            line from CC + (0.5, -dv) to CC + (sx, sy); round;

            linethick = 1.5;
            circle rad 0.42 at CC + (0.2, 0);
            linethick = x;
        B:  CC + (-0.5,  0.0);
        E:  CC + ( 0.5, -d/2);
        C:  CC + ( 0.5,  d/2);
    } )

    ifelse( eval(dir), 1, {
        CC: Q.e  - (0.5,0);
            x = linethick;
            linethick = 2;
            line from CC - (0.025, 0) up_ .20;
            line from CC - (0.025, 0) down_ .20;
            linethick = x;

            line from CC to CC + (-0.5, dv)  then to CC + (-0.5,  d/2);
            line from CC to CC + (-0.5,-dv)  then to CC + (-0.5, -d/2);
            line from CC to CC  + (bx-0.5, 0);

            dr = sqrt((0.5*0.5) + (dv*dv))
            pd = asin(dv/dr);
            dp = 20
            ph =  pd + pi/dp

            sy = 0.25*sin(ph) -dv
            sx = 0.25*cos(ph) - 0.5
            line from CC + (-0.5, -dv) to CC + (sx, sy); round;

            ph = pd - pi/dp
            sy = 0.25*sin(ph) -dv
            sx = 0.25*cos(ph) - 0.5
            line from CC + (-0.5, -dv) to CC + (sx, sy); round;

            linethick = 1.5;
            circle rad 0.42 at CC - (0.2, 0);
            linethick = x;
         B: CC + ( 0.5,  0.0);
         E: CC + (-0.5, -d/2);
         C: CC + (-0.5,  d/2);
    } )
]')

#-----------------------------------------------------------------------
# PNP - bipolarny tranzistor
# bjt_PNP(length_ce, length_b, L|R|U|D)
# length_ce   - dlzka vyvodov medzi C a E
# length_b    - dlzka vyvodu b
# L|R|U|D     - orientacia, todo U|D
#-----------------------------------------------------------------------
define(`bjt_PNP',`[
    ifelse(defn(`d'),  $1, d=1,  d=$1)     # dlzka CE
    ifelse(defn(`bx'), $2, bx=1, bx=$2)    # dlzka bazy
    
    define(dir, index(`RLUP',$3, 0) )    
    Q:box ht d wid 1.5 dotted #invis;
    dx = 0.5;
    dv = 0.3;

    ifelse( eval(dir), 0,       # smer R 
       {
         CC: Q.w  + (0.5,0);
             x = linethick;
            linethick = 2;
            line from CC + (0.025, 0) up_ .20;
            line from CC + (0.025, 0) down_ .20;
            linethick = x;

            line from CC to CC + (0.5, dv)  then to CC + (0.5,  d/2);
            line from CC to CC + (0.5,-dv)  then to CC + (0.5, -d/2);
            line from CC to CC + (0.5-bx, 0);

            dr = sqrt((0.5*0.5) + (dv*dv))
            pd = asin(dv/dr);
            dp = 20
            ph = pi - pd + pi/dp

            sy = 0.25*sin(ph)
            sx = 0.25*cos(ph)
            line from CC to CC + (-sx, sy); round;

            ph = pi - pd - pi/dp
            sy = 0.25*sin(ph)
            sx = 0.25*cos(ph)
            line from CC to CC + (-sx, sy); round;

           linethick = 1.5;
           circle rad 0.42 at CC + (0.2, 0);
           linethick = x;
         B: CC + (-0.5,  0.0);
         C: CC + ( 0.5, -d/2);
         E: CC + ( 0.5,  d/2);
       })

    ifelse( eval(dir), 1,     # smer L
       {
         CC: Q.e  - (0.5,0);
             x = linethick;
        linethick = 2;
        line from CC - (0.025, 0) up_   .20;
        line from CC - (0.025, 0) down_ .20;
        linethick = x;

            line from CC to CC + (-0.5, dv)  then to CC + (-0.5,  d/2);
        line from CC to CC + (-0.5,-dv)  then to CC + (-0.5, -d/2);
            line from CC to CC  + (bx-0.5, 0);

            dr = sqrt((0.5*0.5) + (dv*dv))
            pd = asin(dv/dr);
            dp = 20
        ph =  pd + pi/dp;

            sy = 0.25*sin(ph);
            sx = 0.25*cos(ph);
            line from CC to CC + (-sx, sy); round;

        ph = pd - pi/dp;
            sy = 0.25*sin(ph);
            sx = 0.25*cos(ph);
            line from CC to CC+ (-sx, sy); round;

        linethick = 1.5;
        circle rad 0.42 at CC - (0.2, 0);
        linethick = x;
     B: CC + ( 0.5,  0.0);
     C: CC + (-0.5, -d/2);
         E: CC + (-0.5,  d/2);
       } )
]')



move to 2,2
#test(, A)
right_;
#bjt_PNP(1,1,L)
bjt_NPN(1,1,R)

.PE
