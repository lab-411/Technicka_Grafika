
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(base.ckt)

up_;
I1: source(2,I); llabel(,i_1,);  
    line right_ 1; 
DA: dot; llabel(,a,); line 1;

    move to I1.start; line  right_ 1 ; 
D0: dot; ; 
    line right_ 1; 

    color_red;
    {move to D0; line down_ 0.5; gnd;}
    color_black;

    move to (DA + D0)/2 + (1,0); 
BX: box ht 3 wid 2.5;
    move to (BX.e.x, DA.y); line right_ 1; 
DB: dot; llabel(,b,);

    line -> from DB right_ 1; {"$i_2$" above at last line.c}
    resistor(down_ 2,,E); llabel(,Z,); 
    line left_ 1; 
DG: dot; line to D0;

# popis - sipky
line -> from DA + (0, -0.25) to D0+(0,0.25); "$u_1$" ljust at last line.c;
line -> from DB + (0, -0.25) to DG+(0,0.25); "$u_2$" ljust at last line.c;

.PE
