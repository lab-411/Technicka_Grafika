
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

Origin: Here 
d = 2;

log_init;         # inicializacia makier pre logicke obvody

move to (1,1);
up_; 
H1: Header(2, 6,,,fill_(0.9)); 
"(2,6,,,)" at H1.w rjust;

move to (1,2.5);
H2: Header(1, 6,,,fill_(0.9));
"(1,6,,,)" at H2.w rjust;

move to (1,3.5);
H3: Header(1, 4,0.5,2,fill_(0.9));
"(1,4,0.5,2,)" at H3.w rjust;

move to (4,1.35);
T1: tstrip(R,6,); 
"(R,6)" at T1.e ljust;

move to (4,1.15+1.5);
T2: tstrip(R,6,DO); 
"(R,6,DU)" at T2.e ljust;

move to (4,1.15+2.5);
T2: tstrip(R,4,O; wid=3; ht=.5); 
"(R,4,O;wid=3;ht=.5)" at T2.n above;

"He\\ader()" at (1,0.5);
"ts\\trip()" at (4,0.5);


.PE
