.PS
scale=2.54
cct_init

include(base.ckt)

OA: opamp(,,,,P);
line from OA.V1 up_ .75;
dot;
{line right_ 0.25; capacitor(right_ 1,C+); llabel(,C_1,); rlabel(,10 \mu F,); line .5 then down_ 0.25; gnd;}
line 0.75;
circle rad 0.1; "$V+$" at last circle.n above;

line from OA.V2 down_ .75;
dot;
{line right_ 0.25; reversed(`capacitor', right_, C+); llabel(,C_2,); rlabel(,10 \mu F,); line .5 then down_ 0.25; gnd;}
line 0.75;
circle rad 0.1; "$V-$" at last circle.s below;


.PE
