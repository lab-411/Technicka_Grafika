.PS
scale=2.54
cct_init
include(base.ckt)
B1: box wid 2 ht 2;
line from B1.ne -(0,0.25) right_ 1 ;
P1: circle rad .1; "\textit{P1}" at P1.e ljust;

line from B1.se + (0,0.25) right_ 1 ;
P2: circle rad .1; "\textit{P2}" at P2.e ljust;

"\textit{Output}" at (P1 + P2)/2;

color_red;
"\small{ \"Output\" at (P1 + P2)/2;}" at B1.s + (0,-.2) below ljust;

.PE
