
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


command "\sf"
up_
Orig: Here
move to (Orig+(1,0)); source; { ACsymbol(at last [],,,2:R) }
move to (Orig+(2,0)); source; { DCsymbol(at last [],,,R) }
move to (Orig+(3,0)); battery(,1,R);
move to (Orig+(4,0)); battery(,3,);  rlabel(,,+)

"5V \,\, " at (Orig+(6,0.75)) rjust;  ACsymbol(at last "" ,,,1:R)  
"5V \,\, " at (Orig+(6,1.25)) rjust;  DCsymbol(at last "" ,,,R) 

.PE
