
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_color.ckt)
include(lib_user.ckt)
include(lib_base.ckt)
command"\small \sf"
define(`LF355',`[
    OP: opamp(,,,,);

        line from OP.In1 left_ 0.5;   "2" above ljust;
    INN:last line .end
        line from OP.In2 left_ 0.5;   "3" above ljust;
    INP:last line .end

    P7: 0.25 between OP.N and OP.E;
    P1: 0.5 between OP.N and OP.E;
    P5: 0.75 between OP.N and OP.E;

    P4: 0.5 between OP.S and OP.E;

        line from P7 up_ 0.45; "7" rjust;
    VSP:last line .end;

        line from P4 down_ 0.45; "4" rjust;
    VSN:last line .end;

        line from P1 up_ 0.45; "1" rjust;
    BAL1:last line .end;
        line from P5 up_ 0.45; "5" rjust;
    BAL2:last line .end;
    OUT: OP.Out; "6" at OUT above rjust;
]') 

move to (0,0); 
OP: LF355(); "\sf LF\\355" at OP.OP.se above;
color_red();
#line <- from OP.W left_ 1; ".W" rjust;
line <- from OP.INN left_ 1 up_ .5; ".INN" rjust;
line <- from OP.INP left_ 1 down_ .5; ".INP" rjust;
line <- from OP.VSP up_ 1.25 ; ".VSP" above;
line <- from OP.BAL1 up_ 1 right_ 0.45; ".BAL1" above;
line <- from OP.BAL2 up_ 1 right_ 1.25; ".BAL2" above;
line <- from OP.VSN down_ 0.75 ; ".VSN" below;
line <- from OP.OUT right_ 1; ".OUT" ljust;

move to (6,0); 
right_;
color_black();
OP: LF355();;
box wid (OP.ne-OP.nw).x ht (OP.nw-OP.sw).y at OP.c dashed;
color_blue();
line <- from OP.w left_ 1; ".w" rjust;
line <- from OP.nw left_ 1 up_ 0.5; ".nw" rjust;
line <- from OP.ne right_ 1 up_ 0.5; ".ne" ljust above;
line <- from OP.ne right_ 1 up_ 0.5; ".ne" ljust above;
line <- from OP.se right_ 1 down_ 0.5; ".se" ljust above;
line <- from OP.e right_ 1; ".e" ljust;
line <- from OP.sw left_ 1 down_ 0.5; ".sw" rjust;
line <- from OP.n up_ 1; ".n" above;
line <- from OP.s down_ 1; ".s" below;
line <- from OP.c right_ 0.75 down_ 1.5; ".c" below;

.PE
