
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)
Origin: Here 

d = 2; 
resistor(2,,E); llabel(,R_1,); dot;

linewid = 2.0                      # zmena velkosti komponentu
R1: resistor(3,,ES); llabel(,R_2,); rlabel(,470 \Omega / 5 W,)

dot;                               # zvecseny bod
linewid = 2.54/2                   # uprava rozmerov na standardnu velkost
resistor(d,,E);llabel(,R_3,);      # štandardny rozmer

.PE
