
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


    d = 1.5;

R1: resistor(down_ d,,E); llabel(,R_1,); rarrow(u_{1}, ->, 0.2)
D1: dot; {right_ tconn(,O); "A" ljust;}
R2: resistor(down_ d,,E); llabel(,R_2,); rarrow(u_{2}, ->, 0.2);
D2: dot; {right_ tconn(,O); "B" ljust; }

DC: source(at D1-(2,0)  up_ d); 
   {    DCsymbol(at DC.c,,,R); 
        "$V_0$" at DC.center -(0.6,0); 
        rarrow(u_{0}, <-, 0.3);
    }
    {    line up_ to (Here, R1.start);
         line right_ to R1.start; b_current(i,,,Start, 1.5);
    }
    line from DC.start to (Here, R2.end) then to R2.end;

.PE
