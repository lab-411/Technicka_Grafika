
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


command"\sf"
include(lib_color.ckt)

up_;
move to (0,2);
T: transformer(down_ 2,L,7,W,4);

color_red;
line <- from T.P1 up_ 0.5 left_ 0.5;    ".P1" above rjust;
line <- from T.P2 down_ 0.5 left_ 0.5;  ".P2" below rjust;
line <- from T.S1 up_ 0.5 right_ 0.5;   ".S1" above ljust;
line <- from T.S2 down_ 0.5 right_ 0.5; ".S2" below ljust;
line <- from T.TP left_ 0.75; ".TP"  rjust;
line <- from T.TS right_ 0.75; ".TS"  ljust;

up_;
color_black;
move to (4,2);

T: transformer(down_ 2,L,7,W,4);
color_blue;
B: box wid (T.w-T.e).x ht (T.n-T.s).y at T.c dotted;
line <- from T.sw down_ 0.5 left_ 0.5;   ".sw" below rjust;
line <- from T.nw up_ 0.5 left_ 0.5;     ".nw" above rjust;
line <- from T.ne up_ 0.5 right_ 0.5;    ".ne" above ljust;
line <- from T.se down_ 0.5 right_ 0.5;  ".se" below ljust;
line <- from T.e  right_ 0.75;  ".e" ljust;
line <- from T.w  left_ 0.75;  ".w" rjust;
line <- from T.n  up_ 0.75;  ".n" above;
line <- from T.s  down_ 0.75;  ".s" below;
line <- from T.c  down_ 0.75 right_ 1.25;  ".c" ljust;

.PE
