
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


include(lib_base.ckt)

Origin: Here;             R1: resistor(2,,E);  llabel(,R_1,); "re\\sistor(2,,E)" at R1.start rjust;
move to Origin + (0,1);   C1: capacitor(2);    llabel(,C_1,); "ca\\pacitor(2)" at C1.start rjust;
move to Origin + (0,2);   L1: inductor(2);     llabel(,L_1,); "in\\ductor(2)" at L1.start rjust;
move to Origin + (0,3);   D1: diode(2);        llabel(,D_1,); "di\\ode(2)" at D1.start rjust;

move to Origin + (3,3);   F1: fuse(2);         llabel(,F_1,); "fu\\se(2)" at F1.end ljust;
move to Origin + (3,2);   J1: jumper(2);       llabel(,X_1,); "ju\\mper(2)" at J1.end ljust;
move to Origin + (3,1);   S1: source(2);       "sour\\ce(2)" at S1.end ljust;
move to Origin + (3,0);   B1: battery(2);      "ba\\ttery(2)" at B1.end ljust;

.PE
