
.PS
pi=3.14159265359
                        # parametre z PIC (resp. GNU PIC)
scale = 2.54            # cm - jednotka pre obrazok
maxpswid = 30           # rozmery obrazku
maxpsht = 30            # 30 x 30cm, default je 8.5x11 inch
cct_init                # inicializacia lokalnych premennych

arrowwid  = 0.127       # parametre sipok - sirka
arrowht = 0.254         # dlzka


    right_; 
    resistor(2,,E); llabel(,R_1,); 

    SH:[  
         RR:resistor(2,,ES);
            llabel(,R_2,); rlabel(,470 \Omega / 5 W,);
            box wid elen_ ht elen_*4/5 at RR.center dashed;
        ]
        llabel(,Shield,);  
        { dot(at SH.s); ground;}

        resistor(2,,E); llabel(,R_3,); 

.PE
